library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;

Package constants is
--	constant max_note_cc : natural := 11945;
	constant max_octave : natural := 3;
	constant min_twelfth_cc : natural := 625000;
	constant max_twelfth_cc : natural := 2500000; --2083333
	constant max_note_length_in_twelfths : natural := 96;
	constant max_note_length : natural := max_twelfth_cc * max_note_length_in_twelfths;
	constant sample_rate_cc : natural := 256;
	
	constant num_notes : natural := 12;
	constant music_length : natural := 64;
	constant max_sin_table_index_0 : natural := 1670;
	constant max_sin_table_index_1 : natural := 841;
	constant max_sin_table_index_2 : natural := 425;
	constant max_sin_table_index_3 : natural := 217;
	
	constant note_c : natural := 0;
	constant note_cs : natural := 1;
	constant note_d : natural := 2;
	constant note_ds : natural := 3;
	constant note_e : natural := 4;
	constant note_f : natural := 5;
	constant note_fs : natural := 6;
	constant note_g : natural := 7;
	constant note_gs : natural := 8;
	constant note_a : natural := 9;
	constant note_as : natural := 10;
	constant note_b : natural := 11;
	constant rest : natural := 12;

	type music_pitch_array_type is array(0 to music_length - 1) of unsigned(7 downto 0);
	type music_length_array_type is array(0 to music_length - 1) of unsigned(7 downto 0);
	type sin_table_indices_array_type is array (0 to num_notes + 1) of natural range 0 to max_sin_table_index_0;
	type sin_table_array_type_0 is array (0 to max_sin_table_index_0) of natural range 0 to 255;
	type sin_table_array_type_1 is array (0 to max_sin_table_index_1) of natural range 0 to 255;
	type sin_table_array_type_2 is array (0 to max_sin_table_index_2) of natural range 0 to 255;
	type sin_table_array_type_3 is array (0 to max_sin_table_index_3) of natural range 0 to 255;
	
	signal music_pitch_array : music_pitch_array_type := (x"00", x"02", x"04", x"05", x"07", x"09", x"0B", x"10", x"0B", x"09", x"07", x"05", x"04", x"02", x"00", x"0C", x"10", x"12", x"14", x"15", x"17", x"19", x"1B", x"20", x"1B", x"19", x"17", x"15", x"14", x"12", x"10", x"0C", x"20", x"22", x"24", x"25", x"27", x"29", x"2B", x"30", x"2B", x"29", x"27", x"25", x"24", x"22", x"20", x"0C", x"30", x"32", x"34", x"35", x"37", x"39", x"3B", x"0C", x"3B", x"39", x"37", x"35", x"34", x"32", x"30", x"0C");
	signal music_length_array : music_length_array_type := (x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60");
	constant sin_table_indices_array_0 : sin_table_indices_array_type := (0,187,364,531,688,837,977,1109,1234,1352,1463,1568,1667,1668);
	constant sin_table_indices_array_1 : sin_table_indices_array_type := (0,94,183,267,346,421,491,557,620,679,735,788,838,839);
	constant sin_table_indices_array_2 : sin_table_indices_array_type := (0,47,92,134,174,212,247,280,312,342,370,397,422,423);
	constant sin_table_indices_array_3 : sin_table_indices_array_type := (0,24,47,68,88,107,125,142,158,173,187,201,214,215);
	constant sin_table_array_0 : sin_table_array_type_0 := (0,0,0,0,0,0,1,1,1,1,2,2,3,3,4,4,5,5,6,6,7,8,9,9,10,11,12,13,14,15,16,17,18,19,20,21,23,24,25,27,28,29,31,32,33,35,36,38,39,41,43,44,46,47,49,51,53,54,56,58,60,62,63,65,67,69,71,73,75,77,79,81,83,85,87,89,91,93,95,97,99,101,103,105,108,110,112,114,116,118,120,123,125,127,129,131,133,135,138,140,142,144,146,148,150,152,155,157,159,161,163,165,167,169,171,173,175,177,179,181,183,185,187,189,190,192,194,196,198,200,201,203,205,206,208,210,211,213,215,216,218,219,221,222,224,225,226,228,229,230,232,233,234,235,236,237,238,239,240,241,242,243,244,245,246,247,247,248,249,249,250,251,251,252,252,253,253,253,254,254,254,254,255,255,255,255,255,0,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,7,7,8,9,10,11,12,12,13,14,16,17,18,19,20,21,23,24,25,27,28,30,31,33,34,36,37,39,41,42,44,46,47,49,51,53,55,57,58,60,62,64,66,68,70,72,74,76,79,81,83,85,87,89,91,94,96,98,100,102,105,107,109,111,114,116,118,121,123,125,127,130,132,134,136,139,141,143,145,148,150,152,154,157,159,161,163,165,168,170,172,174,176,178,180,182,184,186,188,190,192,194,196,198,200,202,204,206,207,209,211,213,214,216,217,219,221,222,224,225,227,228,229,231,232,233,235,236,237,238,239,240,241,242,243,244,245,246,247,248,248,249,250,250,251,252,252,252,253,253,254,254,254,254,255,255,255,255,255,0,0,0,0,0,1,1,1,1,2,2,3,3,4,4,5,6,7,7,8,9,10,11,12,13,14,15,16,17,19,20,21,23,24,25,27,28,30,31,33,35,36,38,40,42,43,45,47,49,51,53,55,57,59,61,63,65,67,69,71,74,76,78,80,82,85,87,89,92,94,96,99,101,103,106,108,110,113,115,118,120,122,125,127,130,132,134,137,139,142,144,146,149,151,153,156,158,161,163,165,167,170,172,174,176,179,181,183,185,187,189,192,194,196,198,200,202,204,206,207,209,211,213,215,216,218,220,221,223,225,226,228,229,231,232,233,235,236,237,238,240,241,242,243,244,245,246,247,247,248,249,250,250,251,252,252,253,253,253,254,254,254,255,255,255,255,255,0,0,0,0,0,1,1,1,2,2,3,3,4,4,5,6,6,7,8,9,10,11,12,13,14,16,17,18,20,21,22,24,25,27,28,30,32,33,35,37,39,41,42,44,46,48,50,52,54,57,59,61,63,65,68,70,72,74,77,79,81,84,86,89,91,94,96,98,101,103,106,109,111,114,116,119,121,124,126,129,131,134,137,139,142,144,147,149,152,154,157,159,162,164,167,169,171,174,176,178,181,183,185,188,190,192,194,196,199,201,203,205,207,209,211,213,215,216,218,220,222,223,225,227,228,230,231,233,234,236,237,238,239,241,242,243,244,245,246,247,248,249,249,250,251,251,252,252,253,253,254,254,254,255,255,255,255,0,0,0,0,0,1,1,1,2,2,3,3,4,5,6,6,7,8,9,10,11,12,14,15,16,18,19,20,22,23,25,27,28,30,32,34,35,37,39,41,43,45,47,49,52,54,56,58,61,63,65,68,70,72,75,77,80,82,85,87,90,93,95,98,100,103,106,108,111,114,117,119,122,125,127,130,133,135,138,141,144,146,149,152,154,157,159,162,165,167,170,172,175,177,180,182,185,187,189,192,194,196,199,201,203,205,207,209,212,214,216,217,219,221,223,225,227,228,230,231,233,234,236,237,239,240,241,242,244,245,246,247,248,248,249,250,251,251,252,253,253,254,254,254,255,255,255,255,255,0,0,0,0,1,1,1,2,2,3,3,4,5,5,6,7,8,9,10,11,13,14,15,17,18,20,21,23,24,26,28,30,32,33,35,37,39,42,44,46,48,50,53,55,57,60,62,65,67,70,72,75,78,80,83,86,88,91,94,97,99,102,105,108,111,113,116,119,122,125,128,131,134,136,139,142,145,148,151,153,156,159,162,165,167,170,173,175,178,181,183,186,188,191,193,196,198,200,203,205,207,210,212,214,216,218,220,222,224,226,227,229,231,233,234,236,237,239,240,241,243,244,245,246,247,248,249,250,251,251,252,253,253,254,254,254,255,255,255,255,0,0,0,0,1,1,1,2,2,3,4,4,5,6,7,8,9,10,12,13,14,16,17,19,20,22,24,25,27,29,31,33,35,37,40,42,44,46,49,51,54,56,59,61,64,66,69,72,75,77,80,83,86,89,92,95,97,100,103,106,109,112,115,118,121,125,128,131,134,137,140,143,146,149,152,155,158,161,163,166,169,172,175,178,181,183,186,189,191,194,196,199,202,204,206,209,211,213,216,218,220,222,224,226,228,230,231,233,235,236,238,239,241,242,244,245,246,247,248,249,250,251,251,252,253,253,254,254,254,255,255,255,0,0,0,0,1,1,1,2,3,3,4,5,6,7,8,9,10,12,13,14,16,17,19,21,23,25,26,28,30,33,35,37,39,42,44,47,49,52,54,57,60,62,65,68,71,74,77,80,83,86,89,92,95,98,101,104,107,111,114,117,120,123,127,130,133,136,139,143,146,149,152,155,158,162,165,168,171,174,177,180,183,185,188,191,194,197,199,202,205,207,210,212,214,217,219,221,223,225,227,229,231,233,235,237,238,240,241,243,244,245,246,248,249,250,251,251,252,253,253,254,254,254,255,255,255,0,0,0,0,1,1,2,2,3,4,5,5,6,8,9,10,11,13,14,16,18,20,21,23,25,27,30,32,34,36,39,41,44,46,49,52,55,57,60,63,66,69,72,75,78,82,85,88,91,95,98,101,105,108,111,115,118,121,125,128,132,135,138,142,145,149,152,155,159,162,165,168,172,175,178,181,184,187,190,193,196,199,202,204,207,210,212,215,217,220,222,224,226,228,231,233,234,236,238,240,241,243,244,245,247,248,249,250,251,252,252,253,254,254,254,255,255,255,0,0,0,0,1,1,2,2,3,4,5,6,7,9,10,11,13,14,16,18,20,22,24,26,28,31,33,35,38,41,43,46,49,52,55,58,61,64,67,70,73,77,80,83,87,90,94,97,101,104,108,111,115,119,122,126,129,133,137,140,144,147,151,154,158,161,165,168,172,175,178,182,185,188,191,194,197,200,203,206,209,212,214,217,220,222,224,227,229,231,233,235,237,239,241,242,244,245,246,248,249,250,251,252,253,253,254,254,255,255,255,0,0,0,1,1,1,2,3,4,5,6,7,8,10,11,13,14,16,18,20,22,24,27,29,32,34,37,40,42,45,48,51,54,58,61,64,67,71,74,78,81,85,88,92,96,100,103,107,111,115,118,122,126,130,134,138,141,145,149,153,156,160,164,167,171,175,178,182,185,188,192,195,198,201,205,208,210,213,216,219,221,224,226,229,231,233,235,237,239,241,243,244,246,247,248,250,251,252,252,253,254,254,255,255,255,0,0,0,1,1,2,2,3,4,5,6,8,9,11,12,14,16,18,20,23,25,27,30,33,35,38,41,44,47,50,54,57,60,64,67,71,75,78,82,86,90,94,98,102,106,110,114,118,122,126,130,134,138,142,146,150,154,158,162,166,170,173,177,181,184,188,192,195,198,202,205,208,211,214,217,220,223,225,228,230,233,235,237,239,241,243,244,246,247,249,250,251,252,253,253,254,254,255,255,0,0,0,0);
	constant sin_table_array_1 : sin_table_array_type_1 := (0,0,0,1,1,2,3,4,5,6,7,9,10,12,14,16,18,20,23,25,28,31,33,36,39,43,46,49,53,56,60,63,67,71,75,79,83,87,91,95,99,103,108,112,116,120,125,129,133,138,142,146,150,155,159,163,167,171,175,179,183,187,190,194,198,201,205,208,211,215,218,221,224,226,229,232,234,236,238,240,242,244,246,247,249,250,251,252,253,254,254,255,255,255,0,0,0,1,1,2,3,4,5,7,8,10,12,13,16,18,20,23,25,28,31,34,37,41,44,47,51,55,58,62,66,70,74,79,83,87,91,96,100,105,109,114,118,123,127,132,136,141,145,150,154,159,163,168,172,176,180,184,188,192,196,200,204,207,211,214,217,221,224,227,229,232,235,237,239,241,243,245,247,248,250,251,252,253,254,254,255,255,255,0,0,0,1,1,2,3,4,6,7,9,11,13,15,17,20,23,25,28,31,35,38,42,45,49,53,57,61,65,69,74,78,82,87,92,96,101,106,110,115,120,125,130,134,139,144,149,153,158,163,167,172,176,181,185,189,194,198,202,206,209,213,216,220,223,226,229,232,235,237,240,242,244,246,247,249,250,252,253,253,254,255,255,255,0,0,0,1,2,3,4,5,6,8,10,12,14,17,20,22,25,28,32,35,39,42,46,50,54,59,63,68,72,77,81,86,91,96,101,106,111,116,121,126,131,137,142,147,152,157,162,166,171,176,181,185,190,194,199,203,207,211,215,218,222,225,228,231,234,237,239,242,244,246,248,249,251,252,253,254,254,255,255,0,0,0,1,2,3,4,6,7,9,11,14,16,19,22,25,28,32,35,39,43,47,52,56,61,65,70,75,80,85,90,95,100,106,111,117,122,127,133,138,144,149,154,159,165,170,175,180,185,189,194,199,203,207,212,216,219,223,227,230,233,236,239,241,244,246,248,249,251,252,253,254,255,255,255,0,0,1,1,2,3,5,6,8,10,13,15,18,21,24,28,32,35,39,44,48,53,57,62,67,72,78,83,88,94,99,105,111,116,122,128,134,139,145,151,156,162,167,173,178,183,188,193,198,203,207,212,216,220,224,227,231,234,237,240,243,245,247,249,251,252,253,254,255,255,0,0,1,1,2,4,5,7,9,12,14,17,20,24,27,31,35,40,44,49,54,59,64,69,75,80,86,92,97,103,109,115,121,128,134,140,146,152,158,163,169,175,181,186,191,196,202,206,211,216,220,224,228,231,235,238,241,244,246,248,250,251,253,254,254,255,0,0,1,1,3,4,6,8,10,13,16,19,23,26,30,35,39,44,49,54,60,65,71,77,83,89,95,101,107,114,120,127,133,139,146,152,158,165,171,177,183,188,194,199,205,210,214,219,223,227,231,235,238,241,244,246,249,251,252,253,254,255,255,0,0,1,2,3,5,6,9,11,14,18,21,25,30,34,39,44,49,55,60,66,72,78,85,91,98,105,111,118,125,132,138,145,152,159,165,172,178,184,190,196,202,207,212,217,222,226,231,234,238,241,244,247,249,251,252,254,254,255,0,0,1,2,3,5,7,10,13,16,20,24,28,33,38,43,49,55,61,67,73,80,87,94,101,108,115,122,129,137,144,151,158,165,172,178,185,191,197,203,209,214,220,224,229,233,237,241,244,246,249,251,253,254,255,255,0,0,1,2,4,6,8,11,14,18,22,27,32,37,42,48,54,61,67,74,81,88,96,103,111,118,126,134,141,149,156,164,171,178,185,192,198,205,210,216,221,226,231,235,239,243,246,248,251,252,254,255,255,0,0,1,2,4,6,9,12,16,20,25,30,35,41,47,54,60,67,75,82,90,98,106,114,122,130,138,146,154,162,170,177,184,192,198,205,211,217,223,228,233,237,241,244,247,250,252,253,254,255,0,0,0,0);
	constant sin_table_array_2 : sin_table_array_type_2 := (0,0,1,3,5,7,10,14,18,23,28,33,39,46,53,60,67,75,83,91,99,108,116,125,133,142,150,159,167,175,183,190,198,205,211,218,224,229,234,238,242,246,249,251,253,254,255,0,0,1,3,5,8,12,16,20,25,31,37,44,51,58,66,74,83,91,100,109,118,127,136,145,154,163,172,180,188,196,204,211,217,224,229,235,239,243,247,250,252,254,255,255,0,0,1,3,6,9,13,17,23,28,35,42,49,57,65,74,82,92,101,110,120,130,139,149,158,167,176,185,194,202,209,216,223,229,235,240,244,247,250,253,254,255,0,0,2,4,6,10,14,20,25,32,39,46,54,63,72,81,91,101,111,121,131,142,152,162,171,181,190,199,207,215,222,228,234,239,244,248,251,253,254,255,0,0,2,4,7,11,16,22,28,35,43,52,61,70,80,90,100,111,122,133,144,154,165,175,185,194,203,212,219,227,233,239,244,248,251,253,255,255,0,1,2,5,8,13,18,24,32,39,48,57,67,78,88,99,111,122,134,145,156,167,178,188,198,207,216,224,231,237,243,247,251,253,255,0,1,2,5,9,14,20,27,35,44,54,64,75,86,97,109,121,134,146,158,169,181,191,202,211,220,228,235,241,246,250,253,254,0,1,3,6,10,16,23,30,39,49,60,71,83,95,107,120,133,146,158,171,183,194,205,214,223,231,238,244,249,252,254,255,0,1,3,6,11,18,25,34,44,55,66,78,91,105,118,132,145,159,172,184,196,207,217,226,234,241,247,251,254,255,0,1,3,7,13,20,28,38,49,61,73,87,101,115,129,144,158,172,185,197,209,220,229,237,244,249,253,255,0,1,4,8,14,22,32,42,54,67,81,96,111,126,141,156,171,185,198,210,221,231,239,246,251,254,255,0,1,4,9,16,25,35,47,60,75,90,106,122,138,154,170,184,198,211,223,233,241,247,252,254,0,0,0,0);
	constant sin_table_array_3 : sin_table_array_type_3 := (0,1,5,10,18,28,39,53,67,83,99,116,133,150,167,183,198,211,224,234,242,249,253,255,0,1,5,12,20,31,44,58,74,91,109,127,145,163,180,196,211,224,235,243,250,254,255,0,1,6,13,23,35,49,65,82,101,120,139,158,176,194,209,223,235,244,250,254,0,2,6,14,25,39,54,72,91,111,131,152,171,190,207,222,234,244,251,254,0,2,7,16,28,43,61,80,100,122,144,165,185,203,219,233,244,251,255,0,2,8,18,32,48,67,88,111,134,156,178,198,216,231,243,251,255,0,2,9,20,35,54,75,97,121,146,169,191,211,228,241,250,254,0,3,10,23,39,60,83,107,133,158,183,205,223,238,249,254,0,3,11,25,44,66,91,118,145,172,196,217,234,247,254,0,3,13,28,49,73,101,129,158,185,209,229,244,253,0,4,14,32,54,81,111,141,171,198,221,239,251,255,0,4,16,35,60,90,122,154,184,211,233,247,254,0,0,0,0);
	
end constants;