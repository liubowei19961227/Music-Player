library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity sine_wave_notes is
port( clk: in std_logic;
	  led: out std_logic;
	  s: out std_logic);
end sine_wave_notes;

architecture Behavioral of sine_wave_notes is

constant max_note_cc : integer := 191113;
constant pwm_block_cc : integer := 256;

type note_cc_array_type is array (0 to 11) of integer range 0 to max_note_cc;
type music_array_type is array (0 to 13) of integer range 0 to 11;
type pwm_array_type is array (0 to 11, 0 to 187) of integer range 0 to 255;

constant note_c : integer := 0;
constant note_cs : integer := 1;
constant note_d : integer := 2;
constant note_ds : integer := 3;
constant note_e : integer := 4;
constant note_f : integer := 5;
constant note_fs : integer := 6;
constant note_g : integer := 7;
constant note_gs : integer := 8;
constant note_a : integer := 9;
constant note_as : integer := 10;
constant note_b : integer := 11;

constant note_cc_array : note_cc_array_type := (191113, 180387, 170263, 160707, 151686, 143151, 135137, 127552, 120394, 113636, 107258, 101238);

constant music_array : music_array_type := (note_c, note_d, note_e, note_f, note_g, note_a, note_b, note_c, note_b, note_a, note_g, note_f, note_e, note_d);

constant pwm_array : pwm_array_type := ((0,0,0,0,0,0,1,1,1,1,2,2,3,3,4,4,5,5,6,6,7,8,9,9,10,11,12,13,14,15,16,17,18,19,20,21,23,24,25,26,28,29,30,32,33,35,36,38,39,41,42,44,46,47,49,51,52,54,56,58,59,61,63,65,67,69,71,73,75,76,78,80,82,84,86,88,91,93,95,97,99,101,103,105,107,109,111,114,116,118,120,122,124,126,128,131,133,135,137,139,141,143,145,148,150,152,154,156,158,160,162,164,166,168,170,172,174,176,178,180,182,184,186,188,190,192,193,195,197,199,201,202,204,206,207,209,211,212,214,215,217,218,220,221,223,224,225,227,228,229,231,232,233,234,235,236,237,239,240,241,241,242,243,244,245,246,246,247,248,248,249,250,250,251,251,252,252,252,253,253,253,253,254,254,254,254,254,0),
(0,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,6,7,8,9,10,11,11,12,13,14,16,17,18,19,20,21,23,24,25,27,28,29,31,32,34,36,37,39,40,42,44,45,47,49,51,53,54,56,58,60,62,64,66,68,70,72,74,76,78,80,82,85,87,89,91,93,95,98,100,102,104,107,109,111,113,116,118,120,122,125,127,129,131,134,136,138,140,143,145,147,149,152,154,156,158,160,163,165,167,169,171,173,175,177,180,182,184,186,188,190,192,194,195,197,199,201,203,205,206,208,210,212,213,215,217,218,220,221,223,224,226,227,228,230,231,232,234,235,236,237,238,239,240,241,242,243,244,245,246,247,247,248,249,249,250,251,251,251,252,252,253,253,253,253,254,254,254,254,254,0,0,0,0,0,1,1,1,2,2,2),
(0,0,0,0,0,1,1,1,1,2,2,3,3,4,4,5,6,6,7,8,9,10,11,12,13,14,15,16,17,19,20,21,23,24,25,27,28,30,31,33,35,36,38,40,41,43,45,47,49,51,53,55,57,59,61,63,65,67,69,71,73,75,78,80,82,84,87,89,91,93,96,98,100,103,105,108,110,112,115,117,119,122,124,127,129,131,134,136,139,141,143,146,148,151,153,155,158,160,162,164,167,169,171,174,176,178,180,182,184,187,189,191,193,195,197,199,201,203,205,207,208,210,212,214,216,217,219,221,222,224,225,227,228,230,231,232,234,235,236,238,239,240,241,242,243,244,245,246,247,247,248,249,249,250,251,251,252,252,252,253,253,253,254,254,254,254,254,0,0,0,0,1,1,1,1,2,2,3,3,4,4,5,6,6,7,8,9,10),
(0,0,0,0,0,1,1,1,2,2,3,3,4,4,5,6,6,7,8,9,10,11,12,13,14,16,17,18,19,21,22,24,25,27,28,30,32,33,35,37,39,40,42,44,46,48,50,52,54,56,58,61,63,65,67,70,72,74,76,79,81,83,86,88,91,93,96,98,101,103,106,108,111,113,116,118,121,123,126,128,131,133,136,139,141,144,146,149,151,154,156,159,161,163,166,168,171,173,175,178,180,182,185,187,189,191,193,196,198,200,202,204,206,208,210,212,214,216,217,219,221,223,224,226,227,229,230,232,233,235,236,237,238,240,241,242,243,244,245,246,247,248,248,249,250,250,251,251,252,252,253,253,253,254,254,254,254,0,0,0,0,0,1,1,1,2,2,3,3,4,4,5,6,7,7,8,9,10,11,12,13,14,16,17,18,20,21,22),
(0,0,0,0,0,1,1,1,2,2,3,3,4,5,6,6,7,8,9,10,11,12,14,15,16,17,19,20,22,23,25,26,28,30,32,33,35,37,39,41,43,45,47,49,51,54,56,58,60,63,65,67,70,72,75,77,80,82,85,87,90,92,95,97,100,103,105,108,111,113,116,119,121,124,127,130,132,135,138,140,143,146,148,151,154,156,159,161,164,167,169,172,174,177,179,182,184,186,189,191,193,196,198,200,202,204,207,209,211,213,215,217,219,220,222,224,226,227,229,231,232,234,235,236,238,239,240,241,243,244,245,246,247,248,248,249,250,250,251,252,252,253,253,253,254,254,254,254,254,0,0,0,0,1,1,1,2,2,3,3,4,5,5,6,7,8,9,10,11,12,13,15,16,17,19,20,22,23,25,26,28,30,31,33,35,37,39,41),
(0,0,0,0,1,1,1,2,2,3,3,4,5,5,6,7,8,9,10,11,13,14,15,17,18,20,21,23,24,26,28,30,31,33,35,37,39,41,44,46,48,50,52,55,57,60,62,64,67,70,72,75,77,80,83,85,88,91,93,96,99,102,105,107,110,113,116,119,122,124,127,130,133,136,139,142,144,147,150,153,156,158,161,164,167,169,172,175,177,180,182,185,188,190,192,195,197,200,202,204,207,209,211,213,215,217,219,221,223,225,227,228,230,232,233,235,236,238,239,240,242,243,244,245,246,247,248,249,250,250,251,252,252,253,253,253,254,254,254,254,0,0,0,0,1,1,1,2,2,3,3,4,5,6,6,7,8,9,10,12,13,14,15,17,18,20,21,23,25,26,28,30,32,34,36,38,40,42,44,46,48,51,53,55,58,60,63,65),
(0,0,0,0,1,1,1,2,2,3,4,4,5,6,7,8,9,10,11,13,14,16,17,19,20,22,24,25,27,29,31,33,35,37,39,42,44,46,49,51,53,56,58,61,64,66,69,72,74,77,80,83,85,88,91,94,97,100,103,106,109,112,115,118,121,124,127,130,133,136,139,142,145,148,151,154,157,160,163,166,169,171,174,177,180,183,185,188,191,193,196,198,201,203,206,208,210,212,215,217,219,221,223,225,227,229,230,232,234,235,237,239,240,241,243,244,245,246,247,248,249,250,250,251,252,252,253,253,253,254,254,254,0,0,0,0,1,1,1,2,2,3,4,4,5,6,7,8,9,10,12,13,14,16,17,19,20,22,24,25,27,29,31,33,35,37,39,42,44,46,49,51,53,56,58,61,64,66,69,72,74,77,80,83,86,88,91,94),
(0,0,0,0,1,1,1,2,3,3,4,5,6,7,8,9,10,11,13,14,16,17,19,21,23,24,26,28,30,32,35,37,39,42,44,46,49,51,54,57,59,62,65,68,70,73,76,79,82,85,88,91,94,98,101,104,107,110,113,117,120,123,126,129,133,136,139,142,145,148,152,155,158,161,164,167,170,173,176,179,182,185,188,190,193,196,199,201,204,206,209,211,214,216,218,220,222,225,227,229,230,232,234,236,237,239,240,242,243,244,246,247,248,249,250,250,251,252,252,253,253,253,254,254,254,0,0,0,0,1,1,2,2,3,4,4,5,6,7,8,10,11,12,13,15,17,18,20,22,23,25,27,29,31,33,36,38,40,43,45,47,50,53,55,58,61,63,66,69,72,75,78,81,84,87,90,93,96,99,102,105,108,112,115,118,121,124,127),
(0,0,0,0,1,1,2,2,3,4,5,5,6,8,9,10,11,13,14,16,18,19,21,23,25,27,29,32,34,36,39,41,44,46,49,52,54,57,60,63,66,69,72,75,78,81,84,88,91,94,97,101,104,107,111,114,118,121,124,128,131,135,138,141,145,148,151,155,158,161,164,168,171,174,177,180,183,186,189,192,195,198,201,204,206,209,211,214,216,219,221,223,225,228,230,232,233,235,237,239,240,242,243,244,246,247,248,249,250,251,251,252,253,253,253,254,254,254,0,0,0,1,1,1,2,2,3,4,5,6,7,8,9,11,12,14,15,17,18,20,22,24,26,28,30,33,35,37,40,42,45,47,50,53,56,58,61,64,67,70,73,76,79,83,86,89,92,96,99,102,106,109,112,116,119,122,126,129,133,136,139,143,146,149,153,156,159,163),
(0,0,0,0,1,1,2,2,3,4,5,6,7,9,10,11,13,14,16,18,20,22,24,26,28,31,33,35,38,40,43,46,49,52,54,57,60,64,67,70,73,76,80,83,86,90,93,97,100,104,107,111,114,118,122,125,129,132,136,140,143,147,150,154,157,161,164,168,171,174,178,181,184,187,191,194,197,200,203,205,208,211,214,216,219,221,224,226,228,230,232,234,236,238,240,241,243,244,246,247,248,249,250,251,252,252,253,253,254,254,254,0,0,0,0,1,1,2,3,3,4,5,6,7,9,10,11,13,14,16,18,20,22,24,26,28,31,33,35,38,41,43,46,49,52,55,57,61,64,67,70,73,76,80,83,87,90,93,97,100,104,107,111,115,118,122,125,129,133,136,140,143,147,150,154,157,161,164,168,171,174,178,181,184,188,191,194,197),
(0,0,0,1,1,1,2,3,4,5,6,7,8,10,11,13,14,16,18,20,22,24,27,29,32,34,37,39,42,45,48,51,54,57,61,64,67,70,74,77,81,85,88,92,95,99,103,107,110,114,118,122,126,129,133,137,141,145,148,152,156,159,163,167,170,174,177,181,184,188,191,194,198,201,204,207,210,213,215,218,221,223,226,228,230,232,234,236,238,240,242,243,245,246,247,249,250,251,251,252,253,253,254,254,254,0,0,0,1,1,2,2,3,4,5,6,7,8,10,11,13,15,17,19,21,23,25,27,30,32,35,37,40,43,46,49,52,55,58,61,65,68,71,75,78,82,85,89,93,96,100,104,108,111,115,119,123,127,130,134,138,142,146,149,153,157,160,164,168,171,175,178,182,185,189,192,195,198,201,204,207,210,213,216,219,221,224,226),
(0,0,0,1,1,2,2,3,4,5,6,8,9,11,12,14,16,18,20,22,25,27,30,32,35,38,41,44,47,50,53,57,60,64,67,71,74,78,82,86,90,93,97,101,105,109,113,117,121,125,129,133,137,141,145,149,153,157,161,165,169,173,176,180,184,187,191,194,198,201,204,207,210,213,216,219,222,225,227,230,232,234,236,238,240,242,244,245,247,248,249,250,251,252,252,253,253,254,254,0,0,0,1,1,2,2,3,4,5,7,8,9,11,13,14,16,18,21,23,25,28,30,33,36,38,41,44,47,51,54,57,61,64,68,71,75,79,82,86,90,94,98,102,106,110,114,118,122,126,130,134,138,142,146,150,154,158,162,166,169,173,177,181,184,188,191,195,198,201,205,208,211,214,217,220,222,225,227,230,232,234,236,238,240,242,244,245,247));


constant second_cc : integer := 100000000;

signal pwm_cc : integer range 0 to pwm_block_cc - 1 := 0;
signal pwm_block_partial : integer range 0 to pwm_block_cc - 1 := 0;
signal pwm_block_count : integer range 0 to 192 - 1 := 0;

signal note : integer range 0 to 11 := music_array(0);
signal note_cc : integer range 0 to max_note_cc := pwm_array(note, 0); -- note in clock cycles
signal note_partial : integer range 0 to max_note_cc - 1 := 0;

signal second_partial : integer range 0 to second_cc -1 := 0;
signal second_count : integer range 0 to 13 := 0;

signal square_wave: integer range 0 to 1 := 0;
signal pulse: std_logic := '0';

begin

process (clk)
begin
    if (rising_edge(clk)) then
	     if second_partial = second_cc - 1 then
            second_partial <= 0;
			second_count <= second_count + 1;
			note <= music_array(second_count);
			note_cc <= note_cc_array(note);
			note_partial <= 0;
			square_wave <= 0;
			pwm_block_count <= 0;
			pwm_block_partial <= 0;
			pwm_cc <=  pwm_array(note, 0);
        else
            second_partial <= second_partial + 1;
        end if;
		
		if note_partial = note_cc - 1 then
			note_partial <= 0;
			square_wave <= 1 - square_wave;
			pwm_block_count <= 0;
			pwm_block_partial <= 0;
			pwm_cc <=  pwm_array(note, 0);
			if square_wave = 1 then
				pwm_cc <= pwm_block_cc - pwm_cc;
			end if;
			pulse <= '1';
		else
			note_partial <= note_partial + 1;
        end if;
		
	    if pwm_block_partial = pwm_block_cc - 1 then
            pwm_block_partial <= 0;
			pwm_block_count <= pwm_block_count + 1;
			pwm_cc <=  pwm_array(note, pwm_block_count / 4);
			if square_wave = 1 then
				pwm_cc <= pwm_block_cc - pwm_cc;
			end if;
			pulse <= '1';
        else
            pwm_block_partial <= pwm_block_partial + 1;
		end if;
		
		if pwm_block_partial = pwm_cc then
			pulse <= '0';
		end if;
--		if square_wave = 1 then
--			pulse <= '1';
--		else
--			pulse <= '0';
--		end if;
    end if;
end process;


s <= pulse;
led <= pulse;

end Behavioral;