library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;

Package constants is
--	constant max_note_cc : natural := 11945;
	constant max_octave : natural := 3;
	constant min_twelfth_cc : natural := 500000;
	constant max_twelfth_cc : natural := 3125000; --2083333
	constant max_note_length_in_twelfths : natural := 96;
	constant max_note_length : natural := max_twelfth_cc * max_note_length_in_twelfths;
	constant sample_rate_cc : natural := 256;
	
	constant num_notes : natural := 12;
	constant music_length : natural := 1024;
	constant max_sin_table_index : natural := 3340;
	
	constant note_c : natural := 0;
	constant note_cs : natural := 1;
	constant note_d : natural := 2;
	constant note_ds : natural := 3;
	constant note_e : natural := 4;
	constant note_f : natural := 5;
	constant note_fs : natural := 6;
	constant note_g : natural := 7;
	constant note_gs : natural := 8;
	constant note_a : natural := 9;
	constant note_as : natural := 10;
	constant note_b : natural := 11;
	constant rest : natural := 12;
	
	constant rest_sin_table_index : natural := 3331;

	type music_pitch_array_type is array(0 to music_length - 1) of unsigned(7 downto 0);
	type music_length_array_type is array(0 to music_length - 1) of unsigned(7 downto 0);
	type sin_table_indices_array_type is array (0 to num_notes + 1) of natural range 0 to max_sin_table_index;
	type sin_table_array_type is array (0 to max_sin_table_index) of natural range 0 to 255;
	
	--signal music_pitch_array : music_pitch_array_type := (x"00", x"02", x"04", x"05", x"07", x"09", x"0B", x"10", x"0B", x"09", x"07", x"05", x"04", x"02", x"00", x"0C", x"10", x"12", x"14", x"15", x"17", x"19", x"1B", x"20", x"1B", x"19", x"17", x"15", x"14", x"12", x"10", x"0C", x"20", x"22", x"24", x"25", x"27", x"29", x"2B", x"30", x"2B", x"29", x"27", x"25", x"24", x"22", x"20", x"0C", x"30", x"32", x"34", x"35", x"37", x"39", x"3B", x"0C", x"3B", x"39", x"37", x"35", x"34", x"32", x"30", x"0C");
	--signal music_length_array : music_length_array_type := (x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C");
	constant sin_table_indices_array : sin_table_indices_array_type := (0,374,727,1060,1374,1671,1951,2215,2465,2701,2923,3133,3331,3332);
	constant sin_table_array : sin_table_array_type := (0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,2,2,2,2,2,3,3,3,3,4,4,4,4,5,5,5,5,6,6,6,7,7,8,8,8,9,9,9,10,10,11,11,12,12,12,13,13,14,14,15,15,16,16,17,18,18,19,19,20,20,21,21,22,23,23,24,25,25,26,27,27,28,28,29,30,31,31,32,33,33,34,35,36,36,37,38,39,39,40,41,42,43,43,44,45,46,47,47,48,49,50,51,52,53,53,54,55,56,57,58,59,60,61,62,62,63,64,65,66,67,68,69,70,71,72,73,74,75,76,77,78,79,80,81,82,83,84,85,86,87,88,89,90,91,92,93,94,95,96,97,98,99,100,101,102,103,104,105,107,108,109,110,111,112,113,114,115,116,117,118,119,120,121,123,124,125,126,127,128,129,130,131,132,133,134,135,136,138,139,140,141,142,143,144,145,146,147,148,149,150,151,152,153,155,156,157,158,159,160,161,162,163,164,165,166,167,168,169,170,171,172,173,174,175,176,177,178,179,180,181,182,183,184,185,186,187,188,189,190,190,191,192,193,194,195,196,197,198,199,200,200,201,202,203,204,205,206,206,207,208,209,210,211,211,212,213,214,215,215,216,217,218,218,219,220,221,221,222,223,224,224,225,226,226,227,228,228,229,230,230,231,232,232,233,233,234,235,235,236,236,237,237,238,238,239,239,240,240,241,241,242,242,243,243,244,244,245,245,245,246,246,247,247,247,248,248,248,249,249,249,250,250,250,251,251,251,251,252,252,252,252,253,253,253,253,253,253,254,254,254,254,254,254,254,255,255,255,255,255,255,255,255,255,255,255,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,2,2,2,2,2,3,3,3,3,4,4,4,5,5,5,5,6,6,7,7,7,8,8,8,9,9,10,10,11,11,12,12,12,13,13,14,14,15,16,16,17,17,18,18,19,20,20,21,21,22,23,23,24,25,25,26,27,27,28,29,30,30,31,32,33,33,34,35,36,36,37,38,39,40,41,41,42,43,44,45,46,47,47,48,49,50,51,52,53,54,55,56,57,58,58,59,60,61,62,63,64,65,66,67,68,69,70,71,72,73,74,75,76,78,79,80,81,82,83,84,85,86,87,88,89,90,91,93,94,95,96,97,98,99,100,101,102,104,105,106,107,108,109,110,111,113,114,115,116,117,118,119,121,122,123,124,125,126,127,128,130,131,132,133,134,135,136,138,139,140,141,142,143,144,145,147,148,149,150,151,152,153,154,156,157,158,159,160,161,162,163,164,165,166,168,169,170,171,172,173,174,175,176,177,178,179,180,181,182,183,184,185,186,187,188,189,190,191,192,193,194,195,196,197,198,199,200,201,202,203,204,205,206,206,207,208,209,210,211,212,213,213,214,215,216,217,217,218,219,220,221,221,222,223,224,224,225,226,227,227,228,229,229,230,231,231,232,233,233,234,235,235,236,236,237,238,238,239,239,240,240,241,241,242,242,243,243,244,244,245,245,246,246,246,247,247,248,248,248,249,249,249,250,250,250,251,251,251,252,252,252,252,252,253,253,253,253,253,254,254,254,254,254,254,254,255,255,255,255,255,255,255,255,255,255,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,2,2,2,2,3,3,3,3,4,4,4,4,5,5,5,6,6,7,7,7,8,8,9,9,9,10,10,11,11,12,12,13,13,14,15,15,16,16,17,17,18,19,19,20,21,21,22,23,23,24,25,25,26,27,28,28,29,30,31,31,32,33,34,35,36,36,37,38,39,40,41,42,42,43,44,45,46,47,48,49,50,51,52,53,54,55,56,57,58,59,60,61,62,63,64,65,66,67,68,69,70,71,72,74,75,76,77,78,79,80,81,82,84,85,86,87,88,89,90,92,93,94,95,96,97,99,100,101,102,103,104,106,107,108,109,110,112,113,114,115,116,118,119,120,121,122,124,125,126,127,128,130,131,132,133,134,136,137,138,139,140,142,143,144,145,146,148,149,150,151,152,153,155,156,157,158,159,161,162,163,164,165,166,167,169,170,171,172,173,174,175,176,178,179,180,181,182,183,184,185,186,187,188,189,191,192,193,194,195,196,197,198,199,200,201,202,203,204,205,206,206,207,208,209,210,211,212,213,214,215,216,216,217,218,219,220,221,221,222,223,224,225,225,226,227,228,228,229,230,231,231,232,233,233,234,235,235,236,237,237,238,238,239,240,240,241,241,242,242,243,243,244,244,245,245,246,246,247,247,247,248,248,249,249,249,250,250,250,251,251,251,252,252,252,252,253,253,253,253,253,254,254,254,254,254,254,254,255,255,255,255,255,255,255,255,255,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,2,2,2,2,3,3,3,3,4,4,4,5,5,5,6,6,6,7,7,8,8,9,9,10,10,11,11,12,12,13,13,14,14,15,16,16,17,18,18,19,20,20,21,22,22,23,24,25,25,26,27,28,28,29,30,31,32,33,33,34,35,36,37,38,39,40,41,42,42,43,44,45,46,47,48,49,50,51,52,53,54,56,57,58,59,60,61,62,63,64,65,66,68,69,70,71,72,73,74,76,77,78,79,80,81,83,84,85,86,87,89,90,91,92,94,95,96,97,98,100,101,102,103,105,106,107,109,110,111,112,114,115,116,117,119,120,121,122,124,125,126,128,129,130,131,133,134,135,137,138,139,140,142,143,144,145,147,148,149,150,152,153,154,155,157,158,159,160,162,163,164,165,167,168,169,170,171,173,174,175,176,177,178,180,181,182,183,184,185,186,188,189,190,191,192,193,194,195,196,197,199,200,201,202,203,204,205,206,207,208,209,210,211,212,213,214,215,215,216,217,218,219,220,221,222,223,223,224,225,226,227,227,228,229,230,231,231,232,233,233,234,235,236,236,237,238,238,239,239,240,241,241,242,242,243,243,244,244,245,245,246,246,247,247,248,248,249,249,249,250,250,250,251,251,251,252,252,252,252,253,253,253,253,254,254,254,254,254,254,254,255,255,255,255,255,255,255,255,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,2,2,2,2,3,3,3,3,4,4,4,5,5,6,6,6,7,7,8,8,9,9,10,10,11,11,12,12,13,14,14,15,16,16,17,18,18,19,20,20,21,22,23,23,24,25,26,27,27,28,29,30,31,32,33,34,34,35,36,37,38,39,40,41,42,43,44,45,46,47,48,49,51,52,53,54,55,56,57,58,59,61,62,63,64,65,66,68,69,70,71,72,74,75,76,77,79,80,81,82,84,85,86,87,89,90,91,93,94,95,97,98,99,100,102,103,104,106,107,108,110,111,112,114,115,117,118,119,121,122,123,125,126,127,129,130,131,133,134,135,137,138,139,141,142,144,145,146,148,149,150,152,153,154,155,157,158,159,161,162,163,165,166,167,168,170,171,172,174,175,176,177,179,180,181,182,183,185,186,187,188,189,191,192,193,194,195,196,198,199,200,201,202,203,204,205,206,207,208,209,211,212,213,214,215,216,217,217,218,219,220,221,222,223,224,225,226,227,227,228,229,230,231,231,232,233,234,234,235,236,237,237,238,239,239,240,241,241,242,242,243,244,244,245,245,246,246,247,247,248,248,248,249,249,250,250,250,251,251,251,252,252,252,253,253,253,253,254,254,254,254,254,254,255,255,255,255,255,255,255,255,255,0,0,0,0,0,0,0,0,1,1,1,1,1,1,2,2,2,2,3,3,3,4,4,4,5,5,5,6,6,7,7,8,8,9,9,10,10,11,11,12,13,13,14,15,15,16,17,17,18,19,20,20,21,22,23,24,24,25,26,27,28,29,30,31,32,33,33,34,35,36,37,38,39,41,42,43,44,45,46,47,48,49,50,52,53,54,55,56,57,59,60,61,62,64,65,66,67,69,70,71,72,74,75,76,78,79,80,82,83,84,86,87,88,90,91,92,94,95,97,98,99,101,102,104,105,106,108,109,111,112,113,115,116,118,119,121,122,123,125,126,128,129,131,132,134,135,136,138,139,141,142,144,145,146,148,149,151,152,153,155,156,158,159,160,162,163,165,166,167,169,170,171,173,174,175,177,178,179,181,182,183,184,186,187,188,190,191,192,193,194,196,197,198,199,200,202,203,204,205,206,207,208,210,211,212,213,214,215,216,217,218,219,220,221,222,223,224,225,226,227,227,228,229,230,231,232,233,233,234,235,236,236,237,238,239,239,240,241,241,242,243,243,244,244,245,245,246,247,247,248,248,248,249,249,250,250,251,251,251,252,252,252,253,253,253,253,254,254,254,254,254,254,255,255,255,255,255,255,255,255,0,0,0,0,0,0,0,0,1,1,1,1,1,2,2,2,2,3,3,3,4,4,4,5,5,6,6,7,7,8,8,9,9,10,10,11,12,12,13,13,14,15,16,16,17,18,19,19,20,21,22,23,24,25,25,26,27,28,29,30,31,32,33,34,35,36,37,38,40,41,42,43,44,45,46,48,49,50,51,52,54,55,56,57,59,60,61,62,64,65,66,68,69,70,72,73,75,76,77,79,80,82,83,84,86,87,89,90,92,93,95,96,97,99,100,102,103,105,106,108,109,111,112,114,115,117,118,120,121,123,125,126,128,129,131,132,134,135,137,138,140,141,143,144,146,147,149,150,152,153,155,156,158,159,161,162,163,165,166,168,169,171,172,174,175,176,178,179,181,182,183,185,186,187,189,190,191,193,194,195,196,198,199,200,202,203,204,205,206,208,209,210,211,212,213,214,216,217,218,219,220,221,222,223,224,225,226,227,228,229,230,231,231,232,233,234,235,236,236,237,238,239,239,240,241,242,242,243,244,244,245,245,246,246,247,248,248,249,249,249,250,250,251,251,251,252,252,252,253,253,253,253,254,254,254,254,254,255,255,255,255,255,255,255,0,0,0,0,0,0,0,0,1,1,1,1,1,2,2,2,3,3,3,4,4,4,5,5,6,6,7,7,8,8,9,10,10,11,12,12,13,14,14,15,16,17,17,18,19,20,21,22,23,24,25,25,26,27,28,29,30,32,33,34,35,36,37,38,39,40,42,43,44,45,47,48,49,50,52,53,54,56,57,58,60,61,62,64,65,66,68,69,71,72,74,75,77,78,80,81,83,84,86,87,89,90,92,93,95,96,98,99,101,103,104,106,107,109,111,112,114,115,117,119,120,122,123,125,127,128,130,131,133,135,136,138,139,141,143,144,146,147,149,151,152,154,155,157,158,160,162,163,165,166,168,169,171,172,174,175,177,178,180,181,183,184,185,187,188,190,191,193,194,195,197,198,199,201,202,203,205,206,207,208,210,211,212,213,214,216,217,218,219,220,221,222,223,224,225,226,227,228,229,230,231,232,233,234,235,236,237,237,238,239,240,241,241,242,243,243,244,245,245,246,246,247,248,248,249,249,250,250,251,251,251,252,252,252,253,253,253,254,254,254,254,254,254,255,255,255,255,255,255,255,0,0,0,0,0,0,0,1,1,1,1,1,2,2,2,3,3,3,4,4,5,5,5,6,6,7,8,8,9,9,10,11,11,12,13,14,14,15,16,17,18,19,20,20,21,22,23,24,25,26,27,28,30,31,32,33,34,35,36,38,39,40,41,43,44,45,46,48,49,50,52,53,55,56,57,59,60,62,63,65,66,68,69,71,72,74,75,77,78,80,82,83,85,86,88,90,91,93,95,96,98,100,101,103,105,106,108,110,111,113,115,116,118,120,121,123,125,127,128,130,132,133,135,137,138,140,142,144,145,147,149,150,152,154,155,157,159,160,162,164,165,167,168,170,172,173,175,176,178,179,181,183,184,186,187,189,190,192,193,195,196,197,199,200,202,203,204,206,207,208,210,211,212,214,215,216,217,218,220,221,222,223,224,225,226,227,228,230,231,232,233,233,234,235,236,237,238,239,240,240,241,242,243,243,244,245,245,246,247,247,248,248,249,249,250,250,251,251,252,252,252,253,253,253,254,254,254,254,254,255,255,255,255,255,255,255,0,0,0,0,0,0,0,1,1,1,1,2,2,2,2,3,3,4,4,5,5,6,6,7,7,8,9,9,10,11,11,12,13,14,14,15,16,17,18,19,20,21,22,23,24,25,26,27,28,29,31,32,33,34,35,37,38,39,41,42,43,45,46,47,49,50,52,53,55,56,58,59,61,62,64,65,67,69,70,72,73,75,77,78,80,82,83,85,87,88,90,92,94,95,97,99,101,102,104,106,108,110,111,113,115,117,119,120,122,124,126,128,129,131,133,135,137,138,140,142,144,146,147,149,151,153,154,156,158,160,161,163,165,167,168,170,172,173,175,177,178,180,182,183,185,187,188,190,191,193,194,196,197,199,200,202,203,205,206,208,209,210,212,213,214,216,217,218,220,221,222,223,224,226,227,228,229,230,231,232,233,234,235,236,237,238,239,240,241,241,242,243,244,244,245,246,246,247,248,248,249,249,250,250,251,251,252,252,253,253,253,253,254,254,254,254,255,255,255,255,255,255,0,0,0,0,0,0,1,1,1,1,1,2,2,2,3,3,4,4,5,5,6,6,7,8,8,9,10,10,11,12,13,14,14,15,16,17,18,19,20,21,22,23,24,26,27,28,29,30,32,33,34,36,37,38,40,41,42,44,45,47,48,50,51,53,54,56,58,59,61,62,64,66,67,69,71,72,74,76,78,79,81,83,85,87,88,90,92,94,96,98,100,101,103,105,107,109,111,113,115,117,118,120,122,124,126,128,130,132,134,136,138,139,141,143,145,147,149,151,153,155,156,158,160,162,164,166,167,169,171,173,175,176,178,180,182,183,185,187,188,190,192,193,195,197,198,200,201,203,205,206,208,209,210,212,213,215,216,217,219,220,221,223,224,225,226,228,229,230,231,232,233,234,235,236,237,238,239,240,241,242,243,244,244,245,246,246,247,248,248,249,250,250,251,251,252,252,252,253,253,253,254,254,254,254,255,255,255,255,255,255,0,0,0,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,5,6,6,7,8,8,9,10,11,12,12,13,14,15,16,17,18,19,20,21,23,24,25,26,27,29,30,31,33,34,35,37,38,40,41,43,44,46,47,49,50,52,54,55,57,59,60,62,64,66,67,69,71,73,75,77,78,80,82,84,86,88,90,92,94,96,98,100,102,104,106,108,110,112,114,116,118,120,122,124,126,128,130,132,134,136,138,140,142,144,146,148,150,152,154,156,158,160,162,164,166,168,170,171,173,175,177,179,181,183,184,186,188,190,192,193,195,197,198,200,202,203,205,207,208,210,211,213,214,216,217,219,220,221,223,224,225,227,228,229,230,232,233,234,235,236,237,238,239,240,241,242,243,244,244,245,246,247,247,248,249,249,250,251,251,252,252,252,253,253,253,254,254,254,254,255,255,255,255,255,0,0,0,0,0,0,0,0,0,0);
	
	type twelfth_cc_array_type is array(0 to 255) of integer range 0 to 3200000; 
	constant twelfth_cc_array: twelfth_cc_array_type:=(3125000, 3048780, 2976190, 2906977, 2840909, 2777778, 2717391, 2659574, 2604167, 2551020, 2500000, 2450980, 2403846, 2358491, 2314815, 2272727, 2232143, 2192982, 2155172, 2118644, 2083333, 2049180, 2016129, 1984127, 1953125, 1923077, 1893939, 1865672, 1838235, 1811594, 1785714, 1760563, 1736111, 1712329, 1689189, 1666667, 1644737, 1623377, 1602564, 1582278, 1562500, 1543210, 1524390, 1506024, 1488095, 1470588, 1453488, 1436782, 1420455, 1404494, 1388889, 1373626, 1358696, 1344086, 1329787, 1315789, 1302083, 1288660, 1275510, 1262626, 1250000, 1237624, 1225490, 1213592, 1201923, 1190476, 1179245, 1168224, 1157407, 1146789, 1136364, 1126126, 1116071, 1106195, 1096491, 1086957, 1077586, 1068376, 1059322, 1050420, 1041667, 1033058, 1024590, 1016260, 1008065, 1000000, 992063, 984252, 976563, 968992, 961538, 954198, 946970, 939850, 932836, 925926, 919118, 912409, 905797, 899281, 892857, 886525, 880282, 874126, 868056, 862069, 856164, 850340, 844595, 838926, 833333, 827815, 822368, 816993, 811688, 806452, 801282, 796178, 791139, 786164, 781250, 776398, 771605, 766871, 762195, 757576, 753012, 748503, 744048, 739645, 735294, 730994, 726744, 722543, 718391, 714286, 710227, 706215, 702247, 698324, 694444, 690608, 686813, 683060, 679348, 675676, 672043, 668449, 664894, 661376, 657895, 654450, 651042, 647668, 644330, 641026, 637755, 634518, 631313, 628141, 625000, 621891, 618812, 615764, 612745, 609756, 606796, 603865, 600962, 598086, 595238, 592417, 589623, 586854, 584112, 581395, 578704, 576037, 573394, 570776, 568182, 565611, 563063, 560538, 558036, 555556, 553097, 550661, 548246, 545852, 543478, 541126, 538793, 536481, 534188, 531915, 529661, 527426, 525210, 523013, 520833, 518672, 516529, 514403, 512295, 510204, 508130, 506073, 504032, 502008, 500000, 498008, 496032, 494071, 492126, 490196, 488281, 486381, 484496, 482625, 480769, 478927, 477099, 475285, 473485, 471698, 469925, 468165, 466418, 464684, 462963, 461255, 459559, 457875, 456204, 454545, 452899, 451264, 449640, 448029, 446429, 444840, 443262, 441696, 440141, 438596, 437063, 435540, 434028, 432526, 431034, 429553, 428082, 426621, 425170, 423729);
	
end constants;