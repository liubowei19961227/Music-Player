Package constants is
	constant min_note_cc : natural := 25310;
	constant max_note_cc : natural := 47778;
	constant min_twelfth_cc : natural := 625000;
	constant max_twelfth_cc : natural := 2083333;
end constants;